library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity tb_multiplier_4x4_with_1x1 is
    end tb_multiplier_4x4_with_1x1;
    
    