library ieee;
use ieee.std_logic_1164.all;

entity multiplier_4x4 is
    port (
        
    );
end entity;

architecture structural of multiplier_4x4 is
    
    component multiplier_1x1 is
        port (

        );
    end component multiplier_1x1;
    
    component full_adder is
        port (

        );
    end component full_adder;
    
    signal ;
    begin

end architecture structural;       