library ieee;
use ieee.std_logic_1164.all;

entity multiplier_4x4 is
    port (
        
    );